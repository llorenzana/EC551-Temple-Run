//  ===================================================================================
//  								  Define Module, Inputs and Outputs
//													* 50MHz Clock *
//  ===================================================================================
module ClkDiv_50MHz(
		CLK,
		RST,
		CLKOUT
);

// ====================================================================================
// 										Port Declarations
// ====================================================================================
   input			 CLK;		// 100MHz onboard clock
   input			 RST;		// Reset
   output		 CLKOUT;	// New clock output

// ====================================================================================
// 								Parameters, Register, and Wires
// ====================================================================================
   reg 			 CLKOUT;
	reg 			 flag;

//  ===================================================================================
// 							  				Implementation
//  ===================================================================================

		always @(posedge CLK or posedge RST)
			// Reset clock
			if (RST == 1'b1) 
			begin
				CLKOUT <= 0;
				flag <= 0;
			end
			else 
			begin
				if (flag == 1)
				begin
					CLKOUT <= ~CLKOUT;
					flag <= 0;
				end
				else 
				begin
					flag <= 1;
				end
			end
   
endmodule
