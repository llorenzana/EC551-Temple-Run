`include "intersect_delay.sv"
`include "triangle_intersect.sv"
